    Mac OS X            	   2  �     �                                      ATTR      �   �   �                  �   �  %com.apple.metadata:kMDItemWhereFroms   �     com.apple.provenance   �   <  com.apple.quarantine bplist00�_;https://super-duper-guacamole-q7xvx69x9jwvf9x99.github.dev/_;https://super-duper-guacamole-q7xvx69x9jwvf9x99.github.dev/I                            � �Zx��f�q/0281;695f25b8;Chrome;0A9D3445-7CC9-460A-ACBD-FE09979D085B 
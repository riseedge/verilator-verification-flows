    Mac OS X            	   2  �     �                                      ATTR      �   �   �                  �   �  %com.apple.metadata:kMDItemWhereFroms   �     com.apple.provenance   �   <  com.apple.quarantine bplist00�_;https://super-duper-guacamole-q7xvx69x9jwvf9x99.github.dev/_;https://super-duper-guacamole-q7xvx69x9jwvf9x99.github.dev/I                            � �Zx��f�q/0281;695f25b8;Chrome;F1A78F57-7EF9-465D-BCAE-9A4E0AB3D905 